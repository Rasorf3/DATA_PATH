----------------------------------------------------------------
Library IEEE;
use IEEE.std_logic_1164.all;
----------------------------------------------------------------
entity ALU_n is
generic(
			constant n : natural := 32
			);
port(
		S	 : in std_logic_vector(1 downto 0);
		A,B : in std_logic_vector(n-1 downto 0);
		result : out std_logic_vector(n-1 downto 0)
		);
end entity ALU_n;
----------------------------------------------------------------
architecture struc of ALU_n is
	signal 
begin
	opera_sum : entity work.sumador_n generic map(n) port map(A,B,);
	opera_res : entity work.sumador_n generic map(n) port map(A,B,);
	opera_and : entity work.and_n generic map(n) port map(A,B,);
	opera_or  : entity work.or_n generic map(n) port map(A,B,);
	decode : entity work.mux_4_1x32 port map(S,);
	
end architecture struc;