----------------------------------------------------------
Library IEEE;
use IEEE.std_logic_1164.all;
----------------------------------------------------------
entity decode_1_16 is
port(
		control : in std_logic_vector(4 downto 0);
		D : out std_logic_vector(31 downto 0)
		);
end entity decode_1_16;
----------------------------------------------------------
architecture beh of decode_1_16 is
begin
	process(control) is
		begin
			case(control) is
				
				when "00000" =>
					D<= x"00000001";
				
				when "00001" =>
					D <= x"00000002";
					
				when "00010" =>
					D <= x"00000004";
					
				when "00011" =>
					D <= x"00000008";
					
				when "00100" =>
					D <= x"00000010";
					
				when "00101" =>
					D <= x"00000020";
					
				when "00110" =>
					D <= x"00000040";
					
				when "00111" =>
					D <= x"00000080";
					
				when "01000" =>
					D <= x"00000100";
					
				when "01001" =>
					D <= x"00000200";
					
				when "01010" =>
					D <= x"00000400";
					
				when "01011" =>
					D <= x"00000800";
					
				when "01100" =>
					D <= x"00001000";
					
				when "01101" =>
					D <= x"00002000";
					
				when "01110" =>
					D <= x"00004000";
					
				when "01111" =>
					D <= x"00008000";
					
				when "10000" =>
					D<= x"00010000";
					
				when "10001" =>
					D<= x"00020000";
					
				when "10010" =>
					D<= x"00040000";
					
				when "10011" =>
					D<= x"00080000";
					
				when "10100" =>
					D<= x"00100000";
					
				when "10101" =>
					D<= x"00200000";
					
				when "10110" =>
					D<= x"00400000";
					
				when "10111" =>
					D<= x"00800000";
					
				when "11000" =>
					D<= x"01000000";
					
				when "11001" =>
					D<= x"02000000";
					
				when "11010" =>
					D<= x"04000000";
					
				when "11011" =>
					D<= x"08000000";
					
				when "11100" =>
					D<= x"10000000";
					
				when "11101" =>
					D<= x"20000000";
					
				when "11110" =>
					D<= x"40000000";
					
				when "11111" =>
					D<= x"80000000";
					
									
			end case;
		end process;			
end architecture beh;
----------------------------------------------------------